module DP(start, clk, rst, Vect_E, b_1, b_0, ready,Vect_X, Vect_Y,inc_vector,co);	input start, clk, rst;	output [19:0] Vect_E, b_0, b_1;	output ready, inc_vector;	wire En, inc_counter;	output [19:0] Vect_X, Vect_Y,co;	counter T1 (clk, rst, inc_counter, co);	controller T2 (start, co, clk, rst, En, inc_vector ,inc_counter, ready);	Data_loader T3 (clk, rst, inc_vector, Vect_X, Vect_Y);	Coefficient_calculator T4 (clk, rst, Vect_X, Vect_Y, En, b_0, b_1);	Error_checker T5 (clk, rst, En, Vect_X, Vect_Y, b_1, b_0, Vect_E);endmodule