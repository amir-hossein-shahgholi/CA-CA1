module controller(start, co, clk, rst, En, inc_vector ,inc_counter, ready);	input start, co, clk, rst;	output reg En, inc_vector, inc_counter, ready; 	reg [1:0] ns,ps = 2'b00;	parameter [1:0] Idle=2'b00, Begin=2'b01, Count=2'b10, Ready=2'b11;	always @(ps, start, co) begin		ns=Idle;		ready = 1'b0; inc_counter = 1'b0; inc_vector = 1'b0; En = 1'b0;			case(ps)				Idle: ns= start ? Begin : Idle;				Begin: ns= start ? Begin : Count;				Count: begin ns= co ? Ready : Count; inc_counter= 1'b1; inc_vector = 1'b1; En = 1'b1; end				Ready: begin ns= Ready; ready = 1'b1; end				default:ns = Idle;			endcase	end	always@(posedge clk, posedge rst) begin		if(rst)			ps<=Idle;		else			ps<=ns;	endendmodule